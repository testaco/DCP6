// 2048 x 24 dual-port sine ROM with output registers
// (C) Copyright 2011 John B. Stephensen  All rights reserved.
module Sine2k24 (
   input [10:0] aa,ab,  // address ports
   output [23:0] da,db, // data read ports
   input clk,           // common clock
   input rst            // read port reset
   );
wire [31:0] dal,dam,dah,dbl,dbm,dbh;
// lower block RAM
RAMB16BWER #(
   .DATA_WIDTH_A(9),
   .DATA_WIDTH_B(9),
   .INIT_00(256'hC3AC8E683C09CF904B01B15C02A340D96F008E19A127AA2BAA27A31D97108800),
   .INIT_01(256'h1767A8DAFD131A1400DFB1772FDC7C10991789F14EA0E9275C87AAC3D3DBDBD3),
   .INIT_02(256'hCD770B88F0417EA5B6B39C7030DC74F96BCA1650778C90826333F2A03ECC4AB8),
   .INIT_03(256'hD5C79B52EB68C70A303B29FBB24ECF3580B1C7C4A77121B9389EEB213F45340C),
   .INIT_04(256'hFE1E18EEA02D97DDFFFEDA932A9EF0202E1AE6901982CAF2FAE2AB54DF4A97C5),
   .INIT_05(256'h40686435DB56A7CDC99A42C11641441ECF58B9F203ECAE49BD0B32320DC150BA),
   .INIT_06(256'hFDFCC965CF0811E88F054C62490087DF0903CF6CDB1C2F15CD57B5E6EAC26DEC),
   .INIT_07(256'h47DD3C64540E91DDF2D27BEE2C3407A40D403F0AA002302AF184E5120CD469CC),
   .INIT_08(256'h1CFA9BFF2814C437706C2DB3FD0DE27CDB01EC9D14515520B20A2A11BF357379),
   .INIT_09(256'h9D60E32423E2609E9A57D30F0BC743807E3CBBFBFCBF43889059E4324214A901),
   .INIT_0A(256'h4478671074936D02525E26A9E8E2990C3B27CF345634D0293F12A3F2FEC95198),
   .INIT_0B(256'h112BFC85C5BC6CD2F1C8569D9C53C3EBCC65B8C387053C2CD538552CBD070CCB),
   .INIT_0C(256'hB01024EE6C9E8623747B37A8CFAB3C8380329AB98D17574EFB5E7849D00E03AE),
   .INIT_0D(256'h9B8A2C808741AECEA0265F4BEA3C42FB67875BE21C0BAD030DCA3C623CCB0D04),
   .INIT_0E(256'h34E344571B91B8911B5745E53639EE556E38B5E4C4579C933C98A566D8FDD45E),
   .INIT_0F(256'hD8619C8724727121819357CBF0C64E87700B575503637436A9CEA42B644EE936),
   .INIT_10(256'hE94E642BA4CEA93674630355570B70874EC6F0CB57938121717224879C61D8FF),
   .INIT_11(256'hD4FDD866A5983C939C57C4E4B5386E55EE3936E545571B91B8911B5744E33436),
   .INIT_12(256'h0DCB3C623CCA0D03AD0B1CE25B8767FB423CEA4B5F26A0CEAE4187802C8A9B5E),
   .INIT_13(256'h030ED049785EFB4E57178DB99A3280833CABCFA8377B7423869E6CEE2410B004),
   .INIT_14(256'h0C07BD2C5538D52C3C0587C3B865CCEBC3539C9D56C8F1D26CBCC585FC2B11AE),
   .INIT_15(256'h51C9FEF2A3123F29D0345634CF273B0C99E2E8A9265E52026D937410677844CB),
   .INIT_16(256'hA9144232E459908843BFFCFBBB3C7E8043C70B0FD3579A9E60E22324E3609D98),
   .INIT_17(256'h7335BF112A0AB2205551149DEC01DB7CE20DFDB32D6C7037C41428FF9BFA1C01),
   .INIT_18(256'h69D40C12E584F12A3002A00A3F400DA407342CEE7BD2F2DD910E54643CDD4779),
   .INIT_19(256'h6DC2EAE6B557CD152F1CDB6CCF0309DF870049624C058FE81108CF65C9FCFDCC),
   .INIT_1A(256'h50C10D32320BBD49AEEC03F2B958CF1E444116C1429AC9CDA756DB35646840EC),
   .INIT_1B(256'h974ADF54ABE2FAF2CA821990E61A2E20F09E2A93DAFEFFDD972DA0EE181EFEBA),
   .INIT_1C(256'h34453F21EB9E38B92171A7C4C7B18035CF4EB2FB293B300AC768EB529BC7D5C5),
   .INIT_1D(256'h4ACC3EA0F2336382908C775016CA6BF974DC30709CB3B6A57E41F0880B77CD0C),
   .INIT_1E(256'hDBDBD3C3AA875C27E9A04EF1891799107CDC2F77B1DF00141A13FDDAA86717B8),
   .INIT_1F(256'h8810971DA327AA2BAA27A1198E006FD940A3025CB1014B90CF093C688EACC3D3),
   .INIT_20(256'h3D547298C4F73170B5FF4FA4FE5DC027910072E75FD956D556D95DE369F07800),
   .INIT_21(256'hE999582603EDE6EC00214F89D12484F067E9770FB26017D9A479563D2D25252D),
   .INIT_22(256'h3389F57810BF825B4A4D6490D0248C079536EAB08974707E9DCD0E60C234B648),
   .INIT_23(256'h2B3965AE159839F6D0C5D7054EB231CB804F393C598FDF47C86215DFC1BBCCF4),
   .INIT_24(256'h02E2E81260D369230102266DD66210E0D2E61A70E77E360E061E55AC21B6693B),
   .INIT_25(256'hC0989CCB25AA59333766BE3FEABFBCE231A8470EFD1452B743F5CECEF33FB046),
   .INIT_26(256'h0304379B31F8EF1871FBB49EB7007921F7FD319425E4D1EB33A94B1A163E9314),
   .INIT_27(256'hB923C49CACF26F230E2E8512D4CCF95CF3C0C1F660FED0D60F7C1BEEF42C9734),
   .INIT_28(256'hE4066501D8EC3CC99094D34D03F31E8425FF1463ECAFABE04EF6D6EF41CB8D87),
   .INIT_29(256'h63A01DDCDD1EA06266A92DF1F539BD8082C445050441BD7870A71CCEBEEC57FF),
   .INIT_2A(256'hBC8899F08C6D93FEAEA2DA57181E67F4C5D931CCAACC30D7C1EE5D0E0237AF68),
   .INIT_2B(256'hEFD5047B3B44942E0F38AA6364AD3D15349B483D79FBC4D42BC8ABD443F9F435),
   .INIT_2C(256'h50F0DC1294627ADD8C85C9583155C47D80CE664773E9A9B205A288B730F2FD52),
   .INIT_2D(256'h6576D48079BF523260DAA1B516C4BE059979A51EE4F553FDF336C49EC435F3FC),
   .INIT_2E(256'hCC1DBCA9E56F486FE5A9BB1BCAC712AB92C84B1C3CA9646DC4685B9A28032CA2),
   .INIT_2F(256'h289F6479DC8E8FDF7F6DA935103AB27990F5A9ABFD9D8CCA57325CD59CB217CA),
   .INIT_30(256'h17B29CD55C3257CA8C9DFDABA9F59079B23A1035A96D7FDF8F8EDC79649F2801),
   .INIT_31(256'h2C03289A5B68C46D64A93C1C4BC892AB12C7CA1BBBA9E56F486FE5A9BC1DCCCA),
   .INIT_32(256'hF335C49EC436F3FD53F5E41EA5799905BEC416B5A1DA603252BF7980D47665A2),
   .INIT_33(256'hFDF230B788A205B2A9E9734766CE807DC4553158C9858CDD7A629412DCF050FC),
   .INIT_34(256'hF4F943D4ABC82BD4C4FB793D489B34153DAD6463AA380F2E94443B7B04D5EF52),
   .INIT_35(256'hAF37020E5DEEC1D730CCAACC31D9C5F4671E1857DAA2AEFE936D8CF09988BC35),
   .INIT_36(256'h57ECBECE1CA77078BD41040545C48280BD39F5F12DA96662A01EDDDC1DA06368),
   .INIT_37(256'h8DCB41EFD6F64EE0ABAFEC6314FF25841EF3034DD39490C93CECD8016506E4FF),
   .INIT_38(256'h972CF4EE1B7C0FD6D0FE60F6C1C0F35CF9CCD412852E0E236FF2AC9CC423B987),
   .INIT_39(256'h933E161A4BA933EBD1E4259431FDF7217900B79EB4FB7118EFF8319B37040334),
   .INIT_3A(256'hB03FF3CECEF543B75214FD0E47A831E2BCBFEA3FBE66373359AA25CB9C98C014),
   .INIT_3B(256'h69B621AC551E060E367EE7701AE6D2E01062D66D2602012369D36012E8E20246),
   .INIT_3C(256'hCCBBC1DF1562C847DF8F593C394F80CB31B24E05D7C5D0F6399815AE65392B3B),
   .INIT_3D(256'hB634C2600ECD9D7E707489B0EA3695078C24D090644D4A5B82BF1078F58933F4),
   .INIT_3E(256'h25252D3D5679A4D91760B20F77E967F08424D1894F2100ECE6ED03265899E948),
   .INIT_3F(256'h78F069E35DD956D556D95FE772009127C05DFEA44FFFB57031F7C49872543D2D),
   .DOA_REG(1),
   .DOB_REG(1)
   ) rom0 (
   .ADDRA({aa,3'b000}),
   .DIA(32'h00000000),
   .DIPA(4'h0),
   .DOA(dal),
   .DOPA(),
   .CLKA(clk),
   .WEA(4'h0),
   .ENA(1'b1),
   .REGCEA(1'b1),
   .RSTA(rst),
   .ADDRB({ab,3'b000}),
   .DIB(32'h00000000),
   .DIPB(4'h0),
   .DOB(dbl),
   .DOPB(),
   .CLKB(clk),
   .WEB(4'h0),
   .ENB(1'b1),
   .REGCEB(1'b1),
   .RSTB(rst)
   );
// middle block RAM
RAMB16BWER #(
   .DATA_WIDTH_A(9),
   .DATA_WIDTH_B(9),
   .INIT_00(256'h27C35FFB9733CE6A06A23DD97510AC47E37F1AB651ED8824BF5BF6922DC96400),
   .INIT_01(256'h9633D06D0AA845E27F1BB855F28E2BC864019D39D6720EAB47E37F1BB753EF8B),
   .INIT_02(256'hC76707A645E58423C261009F3EDC7B19B856F59331CF6D0BA947E48220BD5BF8),
   .INIT_03(256'h9E41E48729CC6E11B355F7983ADC7D1FC06102A344E58626C76707A848E88828),
   .INIT_04(256'hFDA54CF29940E68C32D87E24CA6F14BA5F04A84DF2963ADE8226CA6E11B558FB),
   .INIT_05(256'hC97521CD7824CF7A25D07B25D07A24CE7721CA731DC56E17BF6810B86007AF56),
   .INIT_06(256'hE59749FBAC5E0FBF7021D18131E1903FEF9E4CFBA95806B4610FBC6916C3701C),
   .INIT_07(256'h3BF3AC641CD48B42F9B0671DD48A40F5AB6015CA7E33E79B4E02B5691CCE8133),
   .INIT_08(256'hB27131F0B06F2DECAA6826E3A05E1AD793500BC7833EF9B46E29E39D5610C982),
   .INIT_09(256'h35FDC48C5319E0A66C32F7BD82460BCF93571ADDA06326E8AA6C2DEFB07131F2),
   .INIT_0A(256'hB3835323F2C1905F2DFBC9966330FDCA96622DF9C48F5924EEB8814A13DCA56D),
   .INIT_0B(256'h1BF4CCA57D552D04DBB2895F350BE0B58A5F3307DBAF825527FACC9E6F4112E2),
   .INIT_0C(256'h5F422405E7C8A98A6A4A2A09E8C7A68462401DFAD7B4906C4723FED9B38E6841),
   .INIT_0D(256'h76624E39240FF9E3CDB7A089715A422911F8DFC5AC92775D42260BEFD3B69A7D),
   .INIT_0E(256'h584D43382D211509FDF0E3D5C8BAAB9D8E7F6F5F4F3F2E1D0CFAE8D6C3B09D8A),
   .INIT_0F(256'hFFFFFEFDFCFAF8F6F3F0EDE9E5E1DDD8D3CEC8C2BCB5AEA79F978F877E756B62),
   .INIT_10(256'h6B757E878F979FA7AEB5BCC2C8CED3D8DDE1E5E9EDF0F3F6F8FAFCFDFEFFFFFF),
   .INIT_11(256'h9DB0C3D6E8FA0C1D2E3F4F5F6F7F8E9DABBAC8D5E3F0FD0915212D38434D5862),
   .INIT_12(256'h9AB6D3EF0B26425D7792ACC5DFF81129425A7189A0B7CDE3F90F24394E62768A),
   .INIT_13(256'h688EB3D9FE23476C90B4D7FA1D406284A6C7E8092A4A6A8AA9C8E70524425F7D),
   .INIT_14(256'h12416F9ECCFA275582AFDB07335F8AB5E00B355F89B2DB042D557DA5CCF41B41),
   .INIT_15(256'hA5DC134A81B8EE24598FC4F92D6296CAFD306396C9FB2D5F90C1F2235383B3E2),
   .INIT_16(256'h3171B0EF2D6CAAE82663A0DD1A5793CF0B4682BDF7326CA6E019538CC4FD356D),
   .INIT_17(256'hC910569DE3296EB4F93E83C70B5093D71A5EA0E32668AAEC2D6FB0F03171B2F2),
   .INIT_18(256'h81CE1C69B5024E9BE7337ECA1560ABF5408AD41D67B0F9428BD41C64ACF33B82),
   .INIT_19(256'h70C31669BC0F61B40658A9FB4C9EEF3F90E13181D12170BF0F5EACFB4997E533),
   .INIT_1A(256'hAF0760B81068BF176EC51D73CA2177CE247AD0257BD0257ACF2478CD2175C91C),
   .INIT_1B(256'h58B5116ECA2682DE3A96F24DA8045FBA146FCA247ED8328CE64099F24CA5FD56),
   .INIT_1C(256'h88E848A80767C72686E544A30261C01F7DDC3A98F755B3116ECC2987E4419EFB),
   .INIT_1D(256'h5BBD2082E447A90B6DCF3193F556B8197BDC3E9F0061C22384E545A60767C728),
   .INIT_1E(256'hEF53B71B7FE347AB0E72D6399D0164C82B8EF255B81B7FE245A80A6DD03396F8),
   .INIT_1F(256'h64C92D92F65BBF2488ED51B61A7FE347AC1075D93DA2066ACE3397FB5FC3278B),
   .INIT_20(256'hD83CA00468CC3195F95DC2268AEF53B81C81E549AE1277DB40A4096DD2369B00),
   .INIT_21(256'h69CC2F92F557BA1D81E447AA0D71D4379BFE62C6298DF154B81C80E448AC1074),
   .INIT_22(256'h3898F859BA1A7BDC3D9EFF60C12384E647A90A6CCE3092F456B81B7DDF42A407),
   .INIT_23(256'h61BE1B78D63391EE4CAA0867C52382E03F9EFD5CBB1A79D93898F857B71777D7),
   .INIT_24(256'h025AB30D66BF1973CD2781DB3590EB45A0FB57B20D69C5217DD93591EE4AA704),
   .INIT_25(256'h368ADE3287DB3085DA2F84DA2F85DB3188DE358CE23A91E84097EF479FF850A9),
   .INIT_26(256'h1A68B60453A1F0408FDE2E7ECE1F6FC01061B30456A7F94B9EF04396E93C8FE3),
   .INIT_27(256'hC40C539BE32B74BD064F98E22B75BF0A549FEA3581CC1864B1FD4A96E3317ECC),
   .INIT_28(256'h4D8ECE0F4F90D2135597D91C5FA1E5286CAFF4387CC1064B91D61C62A9EF367D),
   .INIT_29(256'hCA023B73ACE61F5993CD08427DB9F4306CA8E5225F9CD9175593D2104F8ECE0D),
   .INIT_2A(256'h4C7CACDC0D3E6FA0D20436699CCF0235699DD2063B70A6DB11477EB5EC235A92),
   .INIT_2B(256'hE40B335A82AAD2FB244D76A0CAF41F4A75A0CCF824507DAAD805336190BEED1D),
   .INIT_2C(256'hA0BDDBFA1837567595B5D5F61738597B9DBFE205284B6F93B8DC01264C7197BE),
   .INIT_2D(256'h899DB1C6DBF0061C32485F768EA5BDD6EE07203A536D88A2BDD9F4102C496582),
   .INIT_2E(256'hA7B2BCC7D2DEEAF6020F1C2A37455462718090A0B0C0D1E2F30517293C4F6275),
   .INIT_2F(256'h00000102030507090C0F12161A1E22272C31373D434A515860687078818A949D),
   .INIT_30(256'h948A817870686058514A433D37312C27221E1A16120F0C090705030201000000),
   .INIT_31(256'h624F3C291705F3E2D1C0B0A0908071625445372A1C0F02F6EADED2C7BCB2A79D),
   .INIT_32(256'h65492C10F4D9BDA2886D533A2007EED6BDA58E765F48321C06F0DBC6B19D8975),
   .INIT_33(256'h97714C2601DCB8936F4B2805E2BF9D7B593817F6D5B59575563718FADBBDA082),
   .INIT_34(256'hEDBE90613305D8AA7D5024F8CCA0754A1FF4CAA0764D24FBD2AA825A330BE4BE),
   .INIT_35(256'h5A23ECB57E4711DBA6703B06D29D693502CF9C693604D2A06F3E0DDCAC7C4C1D),
   .INIT_36(256'hCE8E4F10D2935517D99C5F22E5A86C30F4B97D4208CD93591FE6AC733B02CA92),
   .INIT_37(256'h36EFA9621CD6914B06C17C38F4AF6C28E5A15F1CD9975513D2904F0FCE8E4D0D),
   .INIT_38(256'h7E31E3964AFDB16418CC8135EA9F540ABF752BE2984F06BD742BE39B530CC47D),
   .INIT_39(256'h8F3CE99643F09E4BF9A75604B36110C06F1FCE7E2EDE8F40F0A15304B6681ACC),
   .INIT_3A(256'h50F89F47EF9740E8913AE28C35DE8831DB852FDA842FDA8530DB8732DE8A36E3),
   .INIT_3B(256'hA74AEE9135D97D21C5690DB257FBA045EB9035DB8127CD7319BF660DB35A02A9),
   .INIT_3C(256'h7717B757F89838D9791ABB5CFD9E3FE08223C56708AA4CEE9133D6781BBE6104),
   .INIT_3D(256'hA442DF7D1BB856F49230CE6C0AA947E68423C160FF9E3DDC7B1ABA59F89838D7),
   .INIT_3E(256'h10AC48E4801CB854F18D29C662FE9B37D4710DAA47E4811DBA57F5922FCC6907),
   .INIT_3F(256'h9B36D26D09A440DB7712AE49E5811CB853EF8A26C25DF99531CC6804A03CD874),
   .DOA_REG(1),
   .DOB_REG(1)
   ) rom1 (
   .ADDRA({aa,3'b000}),
   .DIA(32'h00000000),
   .DIPA(4'h0),
   .DOA(dam),
   .DOPA(),
   .CLKA(clk),
   .WEA(4'h0),
   .ENA(1'b1),
   .REGCEA(1'b1),
   .RSTA(rst),
   .ADDRB({ab,3'b000}),
   .DIB(32'h00000000),
   .DIPB(4'h0),
   .DOB(dbm),
   .DOPB(),
   .CLKB(clk),
   .WEB(4'h0),
   .ENB(1'b1),
   .REGCEB(1'b1),
   .RSTB(rst)
   );
// upper block RAM
RAMB16BWER #(
   .DATA_WIDTH_A(9),
   .DATA_WIDTH_B(9),
   .INIT_00(256'h0C0B0B0A0A0A0909090808070707060605050504040303030202010101000000),
   .INIT_01(256'h18181717171616151515141413131312121211111010100F0F0E0E0E0D0D0C0C),
   .INIT_02(256'h242424232322222221212120201F1F1F1E1E1D1D1D1C1C1C1B1B1A1A1A191918),
   .INIT_03(256'h30302F2F2F2E2E2E2D2D2C2C2C2B2B2B2A2A2A29292828282727272626252525),
   .INIT_04(256'h3B3B3B3A3A3A3939393838383737373636363535343434333333323232313130),
   .INIT_05(256'h4646464545454444444343434242424141414040403F3F3F3E3E3E3D3D3D3C3C),
   .INIT_06(256'h5050504F4F4F4F4E4E4E4D4D4D4C4C4C4B4B4B4A4A4A4A494949484848474747),
   .INIT_07(256'h5A59595959585858575757575656565555555554545453535353525252515151),
   .INIT_08(256'h62626261616161606060605F5F5F5F5E5E5E5E5D5D5D5C5C5C5C5B5B5B5B5A5A),
   .INIT_09(256'h6A69696969696868686867676767676666666665656565646464646363636362),
   .INIT_0A(256'h707070706F6F6F6F6F6E6E6E6E6E6D6D6D6D6D6C6C6C6C6C6B6B6B6B6B6A6A6A),
   .INIT_0B(256'h7675757575757575747474747474737373737373727272727271717171717170),
   .INIT_0C(256'h7A7A7A7A79797979797979797878787878787877777777777777767676767676),
   .INIT_0D(256'h7D7D7D7D7D7D7C7C7C7C7C7C7C7C7C7C7C7B7B7B7B7B7B7B7B7B7B7A7A7A7A7A),
   .INIT_0E(256'h7F7F7F7F7F7F7F7F7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7D7D7D7D7D7D7D),
   .INIT_0F(256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F),
   .INIT_10(256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F),
   .INIT_11(256'h7D7D7D7D7D7D7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7F7F7F7F7F7F7F7F7F),
   .INIT_12(256'h7A7A7A7A7B7B7B7B7B7B7B7B7B7B7C7C7C7C7C7C7C7C7C7C7C7D7D7D7D7D7D7D),
   .INIT_13(256'h7676767676777777777777777878787878787879797979797979797A7A7A7A7A),
   .INIT_14(256'h7171717171717272727272737373737373747474747474757575757575757676),
   .INIT_15(256'h6A6A6B6B6B6B6B6C6C6C6C6C6D6D6D6D6D6E6E6E6E6E6F6F6F6F6F7070707070),
   .INIT_16(256'h6363636364646464656565656666666667676767676868686869696969696A6A),
   .INIT_17(256'h5A5B5B5B5B5C5C5C5C5D5D5D5E5E5E5E5F5F5F5F606060606161616162626262),
   .INIT_18(256'h5151525252535353535454545555555556565657575757585858595959595A5A),
   .INIT_19(256'h47474848484949494A4A4A4A4B4B4B4C4C4C4D4D4D4E4E4E4F4F4F4F50505051),
   .INIT_1A(256'h3C3D3D3D3E3E3E3F3F3F40404041414142424243434344444445454546464647),
   .INIT_1B(256'h313132323233333334343435353636363737373838383939393A3A3A3B3B3B3C),
   .INIT_1C(256'h2525262627272728282829292A2A2A2B2B2B2C2C2C2D2D2E2E2E2F2F2F303030),
   .INIT_1D(256'h19191A1A1A1B1B1C1C1C1D1D1D1E1E1F1F1F2020212121222222232324242425),
   .INIT_1E(256'h0C0D0D0E0E0E0F0F101010111112121213131314141515151616171717181818),
   .INIT_1F(256'h000001010102020303030404050505060607070708080909090A0A0A0B0B0C0C),
   .INIT_20(256'hF3F4F4F5F5F5F6F6F6F7F7F8F8F8F9F9FAFAFAFBFBFCFCFCFDFDFEFEFEFFFF00),
   .INIT_21(256'hE7E7E8E8E8E9E9EAEAEAEBEBECECECEDEDEDEEEEEFEFEFF0F0F1F1F1F2F2F3F3),
   .INIT_22(256'hDBDBDBDCDCDDDDDDDEDEDEDFDFE0E0E0E1E1E2E2E2E3E3E3E4E4E5E5E5E6E6E7),
   .INIT_23(256'hCFCFD0D0D0D1D1D1D2D2D3D3D3D4D4D4D5D5D5D6D6D7D7D7D8D8D8D9D9DADADA),
   .INIT_24(256'hC4C4C4C5C5C5C6C6C6C7C7C7C8C8C8C9C9C9CACACBCBCBCCCCCCCDCDCDCECECF),
   .INIT_25(256'hB9B9B9BABABABBBBBBBCBCBCBDBDBDBEBEBEBFBFBFC0C0C0C1C1C1C2C2C2C3C3),
   .INIT_26(256'hAFAFAFB0B0B0B0B1B1B1B2B2B2B3B3B3B4B4B4B5B5B5B5B6B6B6B7B7B7B8B8B8),
   .INIT_27(256'hA5A6A6A6A6A7A7A7A8A8A8A8A9A9A9AAAAAAAAABABABACACACACADADADAEAEAE),
   .INIT_28(256'h9D9D9D9E9E9E9E9F9F9F9FA0A0A0A0A1A1A1A1A2A2A2A3A3A3A3A4A4A4A4A5A5),
   .INIT_29(256'h959696969696979797979898989898999999999A9A9A9A9B9B9B9B9C9C9C9C9D),
   .INIT_2A(256'h8F8F8F8F90909090909191919191929292929293939393939494949494959595),
   .INIT_2B(256'h898A8A8A8A8A8A8A8B8B8B8B8B8B8C8C8C8C8C8C8D8D8D8D8D8E8E8E8E8E8E8F),
   .INIT_2C(256'h8585858586868686868686868787878787878788888888888888898989898989),
   .INIT_2D(256'h8282828282828383838383838383838383848484848484848484848585858585),
   .INIT_2E(256'h8080808080808080818181818181818181818181818181818182828282828282),
   .INIT_2F(256'h8080808080808080808080808080808080808080808080808080808080808080),
   .INIT_30(256'h8080808080808080808080808080808080808080808080808080808080808080),
   .INIT_31(256'h8282828282828181818181818181818181818181818181808080808080808080),
   .INIT_32(256'h8585858584848484848484848484838383838383838383838382828282828282),
   .INIT_33(256'h8989898989888888888888888787878787878786868686868686868585858585),
   .INIT_34(256'h8E8E8E8E8E8E8D8D8D8D8D8C8C8C8C8C8C8B8B8B8B8B8B8A8A8A8A8A8A8A8989),
   .INIT_35(256'h9595949494949493939393939292929292919191919190909090908F8F8F8F8F),
   .INIT_36(256'h9C9C9C9C9B9B9B9B9A9A9A9A9999999998989898989797979796969696969595),
   .INIT_37(256'hA5A4A4A4A4A3A3A3A3A2A2A2A1A1A1A1A0A0A0A09F9F9F9F9E9E9E9E9D9D9D9D),
   .INIT_38(256'hAEAEADADADACACACACABABABAAAAAAAAA9A9A9A8A8A8A8A7A7A7A6A6A6A6A5A5),
   .INIT_39(256'hB8B8B7B7B7B6B6B6B5B5B5B5B4B4B4B3B3B3B2B2B2B1B1B1B0B0B0B0AFAFAFAE),
   .INIT_3A(256'hC3C2C2C2C1C1C1C0C0C0BFBFBFBEBEBEBDBDBDBCBCBCBBBBBBBABABAB9B9B9B8),
   .INIT_3B(256'hCECECDCDCDCCCCCCCBCBCBCACAC9C9C9C8C8C8C7C7C7C6C6C6C5C5C5C4C4C4C3),
   .INIT_3C(256'hDADAD9D9D8D8D8D7D7D7D6D6D5D5D5D4D4D4D3D3D3D2D2D1D1D1D0D0D0CFCFCF),
   .INIT_3D(256'hE6E6E5E5E5E4E4E3E3E3E2E2E2E1E1E0E0E0DFDFDEDEDEDDDDDDDCDCDBDBDBDA),
   .INIT_3E(256'hF3F2F2F1F1F1F0F0EFEFEFEEEEEDEDEDECECECEBEBEAEAEAE9E9E8E8E8E7E7E7),
   .INIT_3F(256'hFFFFFEFEFEFDFDFCFCFCFBFBFAFAFAF9F9F8F8F8F7F7F6F6F6F5F5F5F4F4F3F3),
   .DOA_REG(1),
   .DOB_REG(1)
   ) rom2 (
   .ADDRA({aa,3'b000}),
   .DIA(32'h00000000),
   .DIPA(4'h0),
   .DOA(dah),
   .DOPA(),
   .CLKA(clk),
   .WEA(4'h0),
   .ENA(1'b1),
   .REGCEA(1'b1),
   .RSTA(rst),
   .ADDRB({ab,3'b000}),
   .DIB(32'h00000000),
   .DIPB(4'h0),
   .DOB(dbh),
   .DOPB(),
   .CLKB(clk),
   .WEB(4'h0),
   .ENB(1'b1),
   .REGCEB(1'b1),
   .RSTB(rst)
   );
assign da[7:0] = dal[7:0];
assign da[15:8] = dam[7:0];
assign da[23:16] = dah[7:0];
assign db[7:0] = dbl[7:0];
assign db[15:8] = dbm[7:0];
assign db[23:16] = dbh[7:0];
endmodule
