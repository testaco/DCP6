// 1024 x 18 dual-port half-sine ROM with output registers
// internal RAM output registers not used to minimize delays
// Uses 1 block RAM and 36 registers. 268 MHz maximum clock frequency.
// (C) Copyright 2013 John B. Stephensen  All rights reserved.
module Sine1k2h (
   input [9:0] aa,ab,   // address ports
   output [17:0] da,db, // data read ports
   input clk,           // common clock
   input rst            // read port reset
   );
wire [31:0] dad,dbd;	// RAM data output
wire [3:0] dap,dbp;	// RAM parity output
reg [17:0] qa,qb;		// output registers
// lower block RAM
RAMB16BWER #(
   .DATA_WIDTH_A(18),
   .DATA_WIDTH_B(18),
   .INIT_00(256'h2F1B2BF828D425B1228D1F691C45192115FD12D90FB50C91096D064803240000),
   .INIT_01(256'h613E5E1D5AFC57DB54BA51984E764B544832451041ED3ECB3BA838853562323F),
   .INIT_02(256'h932590098CEC89CF86B2839580777D597A3B771C73FD70DE6DBF6A9F677F645F),
   .INIT_03(256'hC4B1C19BBE85BB6FB858B540B229AF10ABF8A8DFA5C5A2AC9F919C77995C9640),
   .INIT_04(256'hF5C3F2B6EFA8EC9AE98CE67CE36CE05CDD4BDA39D727D415D102CDEECADAC7C6),
   .INIT_05(256'h263E233B20381D341A2F172A1424111D0E150B0D080504FB01F1FEE7FBDBF8D0),
   .INIT_06(256'h5604530D50164D1E4A25472B443141353E393B3D383F354132422F422C412940),
   .INIT_07(256'h84F6820E7F247C3A794F7663737670886D996AA967B964C861D55EE25BEE58F9),
   .INIT_08(256'hB2F9B020AD47AA6CA790A4B4A1D69EF79C17993796559372908F8DAA8AC487DE),
   .INIT_09(256'hDFEFDD28DA60D797D4CDD201CF34CC66C998C6C8C3F6C124BE51BB7DB8A7B5D1),
   .INIT_0A(256'h0BBE090A0655039F00E8FE2FFB75F8BAF5FDF340F081EDC1EB00E83EE57AE2B5),
   .INIT_0B(256'h364933AB310B2E692BC62922267D23D6212E1E841BDA192E168013D211220E70),
   .INIT_0C(256'h5F785CF05A6657DB554E52C050314DA04B0E487A45E5434F40B73E1E3B8338E7),
   .INIT_0D(256'h872F84BF824E7FDB7D667AF0787875FF738471086E8A6C0A698A6707648461FE),
   .INIT_0E(256'hAD58AB01A8A9A650A3F4A1979F399CD99A77981495AF934890E08E768C0B899E),
   .INIT_0F(256'hD1DACF9ECD61CB22C8E2C6A0C45CC216BFCFBD86BB3BB8EFB6A1B451B200AFAC),
   .INIT_10(256'hF49EF27FF05FEE3CEC18E9F2E7CAE5A0E375E148DF19DCE8DAB5D881D64BD413),
   .INIT_11(256'h1590138F118C0F870D810B78096D0761055303430131FF1DFD07FAF0F8D6F6BB),
   .INIT_12(256'h349B32B930D52EEF2D072B1D2931274325542362216E1F791D811B88198D178F),
   .INIT_13(256'h51AC4FEA4E264C604A9848CE47024534436441923FBE3DE83C103A353859367B),
   .INIT_14(256'h6CB16B10696E67C96622647962CE61205F715DC05C0C5A57589F56E5552A536C),
   .INIT_15(256'h8599841B829A81187F937E0C7C837AF7796A77DA764874B4731E71866FEC6E50),
   .INIT_16(256'h9C559AFA999D983D96DB9577941192A8913E8FD18E628CF18B7D8A0788908715),
   .INIT_17(256'hB0D8AFA0AE67AD2BABEDAAADA96AA826A6DFA595A44AA2FCA1ACA05A9F059DAE),
   .INIT_18(256'hC313C201C0ECBFD5BEBBBDA0BC82BB62BA3FB91AB7F3B6C9B59EB470B33FB20D),
   .INIT_19(256'hD2FDD210D120D02FCF3ACE44CD4BCC50CB53CA53C951C84CC746C63CC531C423),
   .INIT_1A(256'hE08ADFC3DEFADE2EDD60DC8FDBBCDAE7DA0FD935D859D77AD699D5B5D4CFD3E7),
   .INIT_1B(256'hEBB4EB13EA70E9CBE923E879E7CCE71DE66CE5B8E502E449E38EE2D1E211E14F),
   .INIT_1C(256'hF472F3F9F37DF2FEF27DF1FAF174F0ECF061EFD4EF44EEB2EE1EED87ECEEEC52),
   .INIT_1D(256'hFAC1FA6EFA19F9C2F968F90CF8ADF84CF7E8F782F719F6AEF641F5D1F55EF4EA),
   .INIT_1E(256'hFE9BFE6FFE42FE12FDDFFDAAFD73FD39FCFCFCBDFC7CFC38FBF2FBA9FB5EFB11),
   .INIT_1F(256'hFFFEFFFAFFF4FFEBFFE0FFD3FFC3FFB0FF9BFF84FF6AFF4DFF2FFF0DFEE9FEC3),
   .INIT_20(256'hFEE9FF0DFF2FFF4DFF6AFF84FF9BFFB0FFC3FFD3FFE0FFEBFFF4FFFAFFFEFFFF),
   .INIT_21(256'hFB5EFBA9FBF2FC38FC7CFCBDFCFCFD39FD73FDAAFDDFFE12FE42FE6FFE9BFEC3),
   .INIT_22(256'hF55EF5D1F641F6AEF719F782F7E8F84CF8ADF90CF968F9C2FA19FA6EFAC1FB11),
   .INIT_23(256'hECEEED87EE1EEEB2EF44EFD4F061F0ECF174F1FAF27DF2FEF37DF3F9F472F4EA),
   .INIT_24(256'hE211E2D1E38EE449E502E5B8E66CE71DE7CCE879E923E9CBEA70EB13EBB4EC52),
   .INIT_25(256'hD4CFD5B5D699D77AD859D935DA0FDAE7DBBCDC8FDD60DE2EDEFADFC3E08AE14F),
   .INIT_26(256'hC531C63CC746C84CC951CA53CB53CC50CD4BCE44CF3AD02FD120D210D2FDD3E7),
   .INIT_27(256'hB33FB470B59EB6C9B7F3B91ABA3FBB62BC82BDA0BEBBBFD5C0ECC201C313C423),
   .INIT_28(256'h9F05A05AA1ACA2FCA44AA595A6DFA826A96AAAADABEDAD2BAE67AFA0B0D8B20D),
   .INIT_29(256'h88908A078B7D8CF18E628FD1913E92A89411957796DB983D999D9AFA9C559DAE),
   .INIT_2A(256'h6FEC7186731E74B4764877DA796A7AF77C837E0C7F938118829A841B85998715),
   .INIT_2B(256'h552A56E5589F5A575C0C5DC05F71612062CE6479662267C9696E6B106CB16E50),
   .INIT_2C(256'h38593A353C103DE83FBE419243644534470248CE4A984C604E264FEA51AC536C),
   .INIT_2D(256'h198D1B881D811F79216E23622554274329312B1D2D072EEF30D532B9349B367B),
   .INIT_2E(256'hF8D6FAF0FD07FF1D0131034305530761096D0B780D810F87118C138F1590178F),
   .INIT_2F(256'hD64BD881DAB5DCE8DF19E148E375E5A0E7CAE9F2EC18EE3CF05FF27FF49EF6BB),
   .INIT_30(256'hB200B451B6A1B8EFBB3BBD86BFCFC216C45CC6A0C8E2CB22CD61CF9ED1DAD413),
   .INIT_31(256'h8C0B8E7690E0934895AF98149A779CD99F39A197A3F4A650A8A9AB01AD58AFAC),
   .INIT_32(256'h64846707698A6C0A6E8A7108738475FF78787AF07D667FDB824E84BF872F899E),
   .INIT_33(256'h3B833E1E40B7434F45E5487A4B0E4DA0503152C0554E57DB5A665CF05F7861FE),
   .INIT_34(256'h112213D21680192E1BDA1E84212E23D6267D29222BC62E69310B33AB364938E7),
   .INIT_35(256'hE57AE83EEB00EDC1F081F340F5FDF8BAFB75FE2F00E8039F0655090A0BBE0E70),
   .INIT_36(256'hB8A7BB7DBE51C124C3F6C6C8C998CC66CF34D201D4CDD797DA60DD28DFEFE2B5),
   .INIT_37(256'h8AC48DAA908F9372965599379C179EF7A1D6A4B4A790AA6CAD47B020B2F9B5D1),
   .INIT_38(256'h5BEE5EE261D564C867B96AA96D99708873767663794F7C3A7F24820E84F687DE),
   .INIT_39(256'h2C412F4232423541383F3B3D3E3941354431472B4A254D1E5016530D560458F9),
   .INIT_3A(256'hFBDBFEE701F104FB08050B0D0E15111D1424172A1A2F1D342038233B263E2940),
   .INIT_3B(256'hCADACDEED102D415D727DA39DD4BE05CE36CE67CE98CEC9AEFA8F2B6F5C3F8D0),
   .INIT_3C(256'h995C9C779F91A2ACA5C5A8DFABF8AF10B229B540B858BB6FBE85C19BC4B1C7C6),
   .INIT_3D(256'h677F6A9F6DBF70DE73FD771C7A3B7D598077839586B289CF8CEC900993259640),
   .INIT_3E(256'h356238853BA83ECB41ED451048324B544E76519854BA57DB5AFC5E1D613E645F),
   .INIT_3F(256'h03240648096D0C910FB512D915FD19211C451F69228D25B128D42BF82F1B323F),
   .INITP_00(256'h5555555555555555555555400000000000000000000000000000000000000000),
   .INITP_01(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9555555555555555555555),
   .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAAAAAAAAA),
   .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
   .INITP_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
   .INITP_05(256'hAAAAAAAAAAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
   .INITP_06(256'h555555555555555555555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
   .INITP_07(256'h0000000000000000000000000000000000000000055555555555555555555555),
   .DOA_REG(0),
   .DOB_REG(0)
   ) rom (
   .ADDRA({aa,4'h0}),
   .DIA(32'h00000000),
   .DIPA(4'h0),
   .DOA(dad),
   .DOPA(dap),
   .CLKA(clk),
   .WEA(4'h0),
   .ENA(1'b1),
   .REGCEA(1'b1),
   .RSTA(rst),
   .ADDRB({ab,4'h0}),
   .DIB(32'h00000000),
   .DIPB(4'h0),
   .DOB(dbd),
   .DOPB(dbp),
   .CLKB(clk),
   .WEB(4'h0),
   .ENB(1'b1),
   .REGCEB(1'b1),
   .RSTB(rst)
   );
// external output registers are faster
always @ (posedge clk)
begin
	qa[15:0] <= dad[15:0];
	qa[17:16] <= dap[1:0];
	qb[15:0] <= dbd[15:0];
	qb[17:16] <= dbp[1:0];
end
// connect outputs
assign da = qa;
assign db = qb;
endmodule
